module bare_processor (
    input logic clk,
    input logic rst,
    input  logic[ 31:0] instruction,
	output logic [31:0] pc_addr,
	output logic [1:0]  im_command,
	input logic [31:0] 	mem2proc_data,
	output logic [31:0] proc2Dmem_addr,
	output logic [1:0] 	proc2Dmem_command,
	output logic [31:0] proc2mem_data,
);

processor proc_module(.clk(clk),
                      .rst(rst),
                      .pipeline_commit_wr_idx(),
                      .pipeline_commit_wr_data(),
                      .pipeline_commit_NPC(),
                      .pipeline_commit_wr(),
                      .instruction(instruction),
                      .pc_addr(pc_addr),
                      .im_command(im_command),
                      .mem2proc_data(mem2proc_data),
                      .proc2Dmem_addr(proc2Dmem_addr),
                      .proc2Dmem_command(proc2Dmem_command),
                      .proc2mem_data(proc2mem_data),
                      .if_PC_out(),
                      .if_NPC_out(),
                      .if_IR_out(),
                      .if_valid_inst_out(),
                      .if_id_PC(),
                      .if_id_NPC(),
                      .if_id_IR(),
                      .if_id_valid_inst(),
                      .id_ex_PC(),
                      .id_ex_NPC(),
                      .id_ex_IR(),
                      .id_ex_valid_inst(),
                      .ex_mem_NPC(),
                      .ex_mem_IR(),
                      .ex_mem_valid_inst(),
                      .mem_wb_NPC(),
                      .mem_wb_IR(),
                      .mem_wb_valid_inst());

endmodule